`ifndef RESOURCES_MUX_SVH
`define RESOURCES_MUX_SVH

import uvm_pkg::*;

package resources_mux;
    //
    `include "uvm_macros.svh"
    `include "./seq_adder_transaction.svh"
    `include "./seq_adder_generator.svh"

endpackage


`endif