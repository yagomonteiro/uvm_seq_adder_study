/*
@author: Yago Monteiro
@brief:  
*/