import uvm_pkg::*;


package ula_resources;
    //
    `include "uvm_macros.svh"
    `include "./ula_agent.svh"
    `include "./ula_driver.svh"
    `include "./ula_env.svh"
    `include "./ula_generator.svh"
    `include "./ula_monitor.svh"
    `include "./ula_scoreboard.svh"
    `include "./ula_transaction.svh"
    `include "./ula_test.sv"      

endpackage


